/* Copyright 2020 pitankar@gmail.com
 * 
 * Permission is hereby granted, free of charge, 
 * to any person obtaining a copy of this software
 * and associated documentation files (the "Software"),
 * to deal in the Software without restriction,
 * including without limitation the rights to use,
 * copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit
 * persons to whom the Software is furnished to do so,
 * subject to the following conditions:
 * 
 * The above copyright notice and this permission
 * notice shall be included in all copies or
 * substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY
 * OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT
 * LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. 
 * IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
 * BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
 * ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE
 * OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 **/

/*
 * Blinks the Green LED on the Lattice ice40 stick
 */
module top(input clk, output g, output r1, r2, r3, r4);
    reg [23:0]   counter;
    reg [0:0]    ff;

    always @(posedge clk) begin
        if (counter == 2000000) 
            begin
            counter <= 0;
            ff[0] <= ~ff[0];
            end
        else 
            counter <= counter + 1;
    end

    assign g = ff[0];
    assign r1 = 1'b0;
    assign r2 = 1'b0;
    assign r3 = 1'b0;
    assign r4 = 1'b0;
endmodule
/* Copyright 2020 pitankar@gmail.com
 * 
 * Permission is hereby granted, free of charge, 
 * to any person obtaining a copy of this software
 * and associated documentation files (the "Software"),
 * to deal in the Software without restriction,
 * including without limitation the rights to use,
 * copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit
 * persons to whom the Software is furnished to do so,
 * subject to the following conditions:
 * 
 * The above copyright notice and this permission
 * notice shall be included in all copies or
 * substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY
 * OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT
 * LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. 
 * IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
 * BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
 * ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE
 * OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 **/

// test bench for transmitter
`timescale 1us/1us

module transmitter_tb;
    reg clk;
    reg [7:0] data;
    wire in_progress;
    reg start;
    wire tx;

    uart_tx transmitter(clk, data, start, in_progress, tx);

    initial begin
        $dumpfile("transmitter_tb.vcd");
        $dumpvars(0,transmitter_tb);

        clk = 1'b0;
        data = 8'b01010101;
        start = 1'b1;
        #20 start = 1'b0;

        #12480 data = 8'b01010101;
        #1248 start = 1'b1;
        #20 start = 1'b0;
        #12480 $finish;
    end

    always begin
        #6 clk = ~clk;
    end
endmodule